27 atime=1442932494.782067
27 ctime=1442932494.787067
